`include "Types.v"

module ID_EXERegister(
    input logic clk,
    input logic rst,
);

endmodule