`include "Types.v"

module ALU();

endmodule