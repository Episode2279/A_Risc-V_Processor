`include "Types.v"

module Extender(
    //not necessary now
);

endmodule