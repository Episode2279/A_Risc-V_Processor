`include "Types.v"

module ExeStages(
    input logic clk,
    input logic rst,
);

endmodule